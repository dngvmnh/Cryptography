
module system (
	clk_clk,
	reset_reset_n,
	led_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[31:0]	led_external_connection_export;
endmodule
